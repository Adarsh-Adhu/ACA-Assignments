`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 25.11.2022 16:42:28
// Design Name: 
// Module Name: MUX_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module MUX16to1_tb();
reg [15:0]i;
reg [3:0]s;
wire f;
MUX16to1 MUX16to1_1(i, s, f);
initial
begin
i=16'b0000000000000001; s=4'b0000; 
#30 i=16'b0000000000000010; s=4'b0001; 
#30 i=16'b0000000000000100; s=4'b0010;
#30 i=16'b0000000000001000; s=4'b0011;
#30 i=16'b0000000000010000; s=4'b0100; 
#30 i=16'b0000000000100000; s=4'b0101; 
#30 i=16'b0000000001000000; s=4'b0110;
#30 i=16'b0000000010000000; s=4'b0111;
#30 i=16'b0000000100000000; s=4'b1000;
#30 i=16'b0000001000000000; s=4'b1001;
#30 i=16'b0000010000000000; s=4'b1010; 
#30 i=16'b0000100000000000; s=4'b1011;
#30 i=16'b0001000000000000; s=4'b1100; 
#30 i=16'b0010000000000000; s=4'b1101; 
#30 i=16'b0100000000000000; s=4'b1110; 
#30 i=16'b1000000000000000; s=4'b1111;
end 
endmodule
